`include "util.svh"

module ir_weights#(
	parameter test_vector_len = 128,
		test_word_width =   16
)(
	output[127: 0][15: 0] weights
);

	//`STATIC_CHECK(test_vector_len == 128, "Invalid vector length, expected: 128");
	//`STATIC_CHECK(test_word_width == 16, "Invalid word length, expected: 16");

	assign weights[0] = 16'h05C2;
	assign weights[1] = 16'h0B8D;
	assign weights[2] = 16'h0E84;
	assign weights[3] = 16'h105B;
	assign weights[4] = 16'h0EF7;
	assign weights[5] = 16'h09DD;
	assign weights[6] = 16'h04A1;
	assign weights[7] = 16'hFF3F;
	assign weights[8] = 16'hFA52;
	assign weights[9] = 16'hF83B;
	assign weights[10] = 16'hF89C;
	assign weights[11] = 16'hFB69;
	assign weights[12] = 16'hFEFA;
	assign weights[13] = 16'h02A5;
	assign weights[14] = 16'h058B;
	assign weights[15] = 16'h07DD;
	assign weights[16] = 16'h07EC;
	assign weights[17] = 16'h0640;
	assign weights[18] = 16'h04A6;
	assign weights[19] = 16'h02B5;
	assign weights[20] = 16'hFFE4;
	assign weights[21] = 16'hFF51;
	assign weights[22] = 16'hFF28;
	assign weights[23] = 16'hFEA7;
	assign weights[24] = 16'hFFCC;
	assign weights[25] = 16'h0107;
	assign weights[26] = 16'h0173;
	assign weights[27] = 16'h01A9;
	assign weights[28] = 16'h01A8;
	assign weights[29] = 16'h0119;
	assign weights[30] = 16'h00B1;
	assign weights[31] = 16'hFFD2;
	assign weights[32] = 16'hFE9D;
	assign weights[33] = 16'hFDC4;
	assign weights[34] = 16'hFD29;
	assign weights[35] = 16'hFCB9;
	assign weights[36] = 16'hFCAF;
	assign weights[37] = 16'hFCC7;
	assign weights[38] = 16'hFC88;
	assign weights[39] = 16'hFCC3;
	assign weights[40] = 16'hFD7E;
	assign weights[41] = 16'hFE02;
	assign weights[42] = 16'hFEA8;
	assign weights[43] = 16'hFF97;
	assign weights[44] = 16'h0086;
	assign weights[45] = 16'h00B9;
	assign weights[46] = 16'h00B0;
	assign weights[47] = 16'h0083;
	assign weights[48] = 16'h0028;
	assign weights[49] = 16'h0042;
	assign weights[50] = 16'h000D;
	assign weights[51] = 16'hFFA3;
	assign weights[52] = 16'hFFA2;
	assign weights[53] = 16'hFF36;
	assign weights[54] = 16'hFE60;
	assign weights[55] = 16'hFDE1;
	assign weights[56] = 16'hFDBA;
	assign weights[57] = 16'hFDE6;
	assign weights[58] = 16'hFE49;
	assign weights[59] = 16'hFF1E;
	assign weights[60] = 16'h0028;
	assign weights[61] = 16'h010E;
	assign weights[62] = 16'h01F1;
	assign weights[63] = 16'h021C;
	assign weights[64] = 16'h01A7;
	assign weights[65] = 16'h0085;
	assign weights[66] = 16'hFF10;
	assign weights[67] = 16'hFDE7;
	assign weights[68] = 16'hFD23;
	assign weights[69] = 16'hFCEF;
	assign weights[70] = 16'hFD11;
	assign weights[71] = 16'hFD44;
	assign weights[72] = 16'hFDAB;
	assign weights[73] = 16'hFE18;
	assign weights[74] = 16'hFE3C;
	assign weights[75] = 16'hFE26;
	assign weights[76] = 16'hFE18;
	assign weights[77] = 16'hFE30;
	assign weights[78] = 16'hFE6E;
	assign weights[79] = 16'hFECD;
	assign weights[80] = 16'hFF55;
	assign weights[81] = 16'hFFB9;
	assign weights[82] = 16'hFFEA;
	assign weights[83] = 16'h001D;
	assign weights[84] = 16'h0015;
	assign weights[85] = 16'hFFBF;
	assign weights[86] = 16'hFF77;
	assign weights[87] = 16'hFF36;
	assign weights[88] = 16'hFEF0;
	assign weights[89] = 16'hFEE1;
	assign weights[90] = 16'hFEAA;
	assign weights[91] = 16'hFE68;
	assign weights[92] = 16'hFE3A;
	assign weights[93] = 16'hFE45;
	assign weights[94] = 16'hFE28;
	assign weights[95] = 16'hFE06;
	assign weights[96] = 16'hFE10;
	assign weights[97] = 16'hFE4C;
	assign weights[98] = 16'hFEA4;
	assign weights[99] = 16'hFEE8;
	assign weights[100] = 16'hFEFF;
	assign weights[101] = 16'hFF05;
	assign weights[102] = 16'hFF0A;
	assign weights[103] = 16'hFF00;
	assign weights[104] = 16'hFF06;
	assign weights[105] = 16'hFF06;
	assign weights[106] = 16'hFEFA;
	assign weights[107] = 16'hFEE6;
	assign weights[108] = 16'hFEBD;
	assign weights[109] = 16'hFE66;
	assign weights[110] = 16'hFDE8;
	assign weights[111] = 16'hFD85;
	assign weights[112] = 16'hFD60;
	assign weights[113] = 16'hFD97;
	assign weights[114] = 16'hFE17;
	assign weights[115] = 16'hFEBA;
	assign weights[116] = 16'hFF3C;
	assign weights[117] = 16'hFF8B;
	assign weights[118] = 16'hFF90;
	assign weights[119] = 16'hFF5C;
	assign weights[120] = 16'hFF17;
	assign weights[121] = 16'hFED0;
	assign weights[122] = 16'hFE7E;
	assign weights[123] = 16'hFE31;
	assign weights[124] = 16'hFDF9;
	assign weights[125] = 16'hFDD7;
	assign weights[126] = 16'hFDD9;
	assign weights[127] = 16'hFDFD;
endmodule
