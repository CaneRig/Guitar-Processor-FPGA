module ir_weights(
     output[255: 0][15: 0] weights;
);
	assign weights[0] = 16'h0519;
	assign weights[1] = 16'h0B13;
	assign weights[2] = 16'h0E31;
	assign weights[3] = 16'h1021;
	assign weights[4] = 16'h0ECA;
	assign weights[5] = 16'h09AD;
	assign weights[6] = 16'h0468;
	assign weights[7] = 16'hFF08;
	assign weights[8] = 16'hFA23;
	assign weights[9] = 16'hF818;
	assign weights[10] = 16'hF880;
	assign weights[11] = 16'hFB49;
	assign weights[12] = 16'hFECD;
	assign weights[13] = 16'h0264;
	assign weights[14] = 16'h053B;
	assign weights[15] = 16'h0781;
	assign weights[16] = 16'h0782;
	assign weights[17] = 16'h05C5;
	assign weights[18] = 16'h0422;
	assign weights[19] = 16'h023A;
	assign weights[20] = 16'hFF85;
	assign weights[21] = 16'hFF0A;
	assign weights[22] = 16'hFEF3;
	assign weights[23] = 16'hFE78;
	assign weights[24] = 16'hFF91;
	assign weights[25] = 16'h00BC;
	assign weights[26] = 16'h011D;
	assign weights[27] = 16'h0154;
	assign weights[28] = 16'h0163;
	assign weights[29] = 16'h00F7;
	assign weights[30] = 16'h00B9;
	assign weights[31] = 16'hFFF3;
	assign weights[32] = 16'hFEC6;
	assign weights[33] = 16'hFDF9;
	assign weights[34] = 16'hFD60;
	assign weights[35] = 16'hFCE0;
	assign weights[36] = 16'hFCCF;
	assign weights[37] = 16'hFCF2;
	assign weights[38] = 16'hFCBC;
	assign weights[39] = 16'hFCF2;
	assign weights[40] = 16'hFDA5;
	assign weights[41] = 16'hFE1B;
	assign weights[42] = 16'hFEA8;
	assign weights[43] = 16'hFF77;
	assign weights[44] = 16'h004A;
	assign weights[45] = 16'h0071;
	assign weights[46] = 16'h006C;
	assign weights[47] = 16'h0043;
	assign weights[48] = 16'hFFEB;
	assign weights[49] = 16'hFFFC;
	assign weights[50] = 16'hFFB7;
	assign weights[51] = 16'hFF40;
	assign weights[52] = 16'hFF3B;
	assign weights[53] = 16'hFECD;
	assign weights[54] = 16'hFDEF;
	assign weights[55] = 16'hFD67;
	assign weights[56] = 16'hFD3C;
	assign weights[57] = 16'hFD67;
	assign weights[58] = 16'hFDC6;
	assign weights[59] = 16'hFE87;
	assign weights[60] = 16'hFF70;
	assign weights[61] = 16'h0036;
	assign weights[62] = 16'h0101;
	assign weights[63] = 16'h0116;
	assign weights[64] = 16'h0090;
	assign weights[65] = 16'hFF6B;
	assign weights[66] = 16'hFE0B;
	assign weights[67] = 16'hFD0D;
	assign weights[68] = 16'hFC8C;
	assign weights[69] = 16'hFCA3;
	assign weights[70] = 16'hFD06;
	assign weights[71] = 16'hFD67;
	assign weights[72] = 16'hFDDA;
	assign weights[73] = 16'hFE47;
	assign weights[74] = 16'hFE64;
	assign weights[75] = 16'hFE2A;
	assign weights[76] = 16'hFDED;
	assign weights[77] = 16'hFDED;
	assign weights[78] = 16'hFE29;
	assign weights[79] = 16'hFE8C;
	assign weights[80] = 16'hFF1E;
	assign weights[81] = 16'hFF84;
	assign weights[82] = 16'hFFA3;
	assign weights[83] = 16'hFFB8;
	assign weights[84] = 16'hFF9A;
	assign weights[85] = 16'hFF38;
	assign weights[86] = 16'hFEED;
	assign weights[87] = 16'hFEC2;
	assign weights[88] = 16'hFEA1;
	assign weights[89] = 16'hFEBA;
	assign weights[90] = 16'hFE9B;
	assign weights[91] = 16'hFE55;
	assign weights[92] = 16'hFE13;
	assign weights[93] = 16'hFE0A;
	assign weights[94] = 16'hFDDE;
	assign weights[95] = 16'hFDB9;
	assign weights[96] = 16'hFDDA;
	assign weights[97] = 16'hFE3A;
	assign weights[98] = 16'hFEB7;
	assign weights[99] = 16'hFF18;
	assign weights[100] = 16'hFF39;
	assign weights[101] = 16'hFF3A;
	assign weights[102] = 16'hFF31;
	assign weights[103] = 16'hFF14;
	assign weights[104] = 16'hFF02;
	assign weights[105] = 16'hFEF3;
	assign weights[106] = 16'hFEEE;
	assign weights[107] = 16'hFEE6;
	assign weights[108] = 16'hFEC2;
	assign weights[109] = 16'hFE7A;
	assign weights[110] = 16'hFE17;
	assign weights[111] = 16'hFDD3;
	assign weights[112] = 16'hFDCB;
	assign weights[113] = 16'hFE18;
	assign weights[114] = 16'hFEAA;
	assign weights[115] = 16'hFF5F;
	assign weights[116] = 16'hFFF9;
	assign weights[117] = 16'h005E;
	assign weights[118] = 16'h0074;
	assign weights[119] = 16'h0045;
	assign weights[120] = 16'hFFFE;
	assign weights[121] = 16'hFFAE;
	assign weights[122] = 16'hFF46;
	assign weights[123] = 16'hFEDF;
	assign weights[124] = 16'hFE94;
	assign weights[125] = 16'hFE63;
	assign weights[126] = 16'hFE51;
	assign weights[127] = 16'hFE6B;
	assign weights[128] = 16'hFEB9;
	assign weights[129] = 16'hFF17;
	assign weights[130] = 16'hFF6A;
	assign weights[131] = 16'hFF9B;
	assign weights[132] = 16'hFFCD;
	assign weights[133] = 16'h0006;
	assign weights[134] = 16'h003C;
	assign weights[135] = 16'h008E;
	assign weights[136] = 16'h0102;
	assign weights[137] = 16'h0149;
	assign weights[138] = 16'h0161;
	assign weights[139] = 16'h0140;
	assign weights[140] = 16'h00C9;
	assign weights[141] = 16'h003C;
	assign weights[142] = 16'hFFAE;
	assign weights[143] = 16'hFF44;
	assign weights[144] = 16'hFF24;
	assign weights[145] = 16'hFF39;
	assign weights[146] = 16'hFF59;
	assign weights[147] = 16'hFF79;
	assign weights[148] = 16'hFF6F;
	assign weights[149] = 16'hFF4E;
	assign weights[150] = 16'hFF23;
	assign weights[151] = 16'hFF03;
	assign weights[152] = 16'hFF0D;
	assign weights[153] = 16'hFF36;
	assign weights[154] = 16'hFF69;
	assign weights[155] = 16'hFF8E;
	assign weights[156] = 16'hFF98;
	assign weights[157] = 16'hFF7A;
	assign weights[158] = 16'hFF43;
	assign weights[159] = 16'hFF1D;
	assign weights[160] = 16'hFF0C;
	assign weights[161] = 16'hFF05;
	assign weights[162] = 16'hFF2A;
	assign weights[163] = 16'hFF6D;
	assign weights[164] = 16'hFFC1;
	assign weights[165] = 16'h000B;
	assign weights[166] = 16'h002B;
	assign weights[167] = 16'h0025;
	assign weights[168] = 16'hFFF3;
	assign weights[169] = 16'hFF92;
	assign weights[170] = 16'hFF30;
	assign weights[171] = 16'hFEFA;
	assign weights[172] = 16'hFEEB;
	assign weights[173] = 16'hFF13;
	assign weights[174] = 16'hFF65;
	assign weights[175] = 16'hFFB7;
	assign weights[176] = 16'h0007;
	assign weights[177] = 16'h0059;
	assign weights[178] = 16'h0097;
	assign weights[179] = 16'h00AD;
	assign weights[180] = 16'h00B1;
	assign weights[181] = 16'h00B6;
	assign weights[182] = 16'h00BA;
	assign weights[183] = 16'h009F;
	assign weights[184] = 16'h0069;
	assign weights[185] = 16'h0024;
	assign weights[186] = 16'hFFD7;
	assign weights[187] = 16'hFF95;
	assign weights[188] = 16'hFF69;
	assign weights[189] = 16'hFF6A;
	assign weights[190] = 16'hFF9D;
	assign weights[191] = 16'hFFEF;
	assign weights[192] = 16'h0056;
	assign weights[193] = 16'h00BB;
	assign weights[194] = 16'h0107;
	assign weights[195] = 16'h0141;
	assign weights[196] = 16'h0153;
	assign weights[197] = 16'h013F;
	assign weights[198] = 16'h011D;
	assign weights[199] = 16'h00F9;
	assign weights[200] = 16'h00EA;
	assign weights[201] = 16'h00E8;
	assign weights[202] = 16'h00E7;
	assign weights[203] = 16'h00EC;
	assign weights[204] = 16'h00F1;
	assign weights[205] = 16'h00FC;
	assign weights[206] = 16'h0105;
	assign weights[207] = 16'h00F8;
	assign weights[208] = 16'h00DC;
	assign weights[209] = 16'h00C9;
	assign weights[210] = 16'h00B9;
	assign weights[211] = 16'h0092;
	assign weights[212] = 16'h0065;
	assign weights[213] = 16'h0047;
	assign weights[214] = 16'h002F;
	assign weights[215] = 16'h0023;
	assign weights[216] = 16'h0029;
	assign weights[217] = 16'h0031;
	assign weights[218] = 16'h0033;
	assign weights[219] = 16'h0043;
	assign weights[220] = 16'h0061;
	assign weights[221] = 16'h0079;
	assign weights[222] = 16'h0080;
	assign weights[223] = 16'h0080;
	assign weights[224] = 16'h0073;
	assign weights[225] = 16'h005C;
	assign weights[226] = 16'h0046;
	assign weights[227] = 16'h0035;
	assign weights[228] = 16'h0038;
	assign weights[229] = 16'h0043;
	assign weights[230] = 16'h0052;
	assign weights[231] = 16'h0066;
	assign weights[232] = 16'h007C;
	assign weights[233] = 16'h007E;
	assign weights[234] = 16'h006F;
	assign weights[235] = 16'h0058;
	assign weights[236] = 16'h004A;
	assign weights[237] = 16'h0045;
	assign weights[238] = 16'h004C;
	assign weights[239] = 16'h0059;
	assign weights[240] = 16'h005E;
	assign weights[241] = 16'h005A;
	assign weights[242] = 16'h0051;
	assign weights[243] = 16'h0037;
	assign weights[244] = 16'h0005;
	assign weights[245] = 16'hFFC7;
	assign weights[246] = 16'hFF8B;
	assign weights[247] = 16'hFF5D;
	assign weights[248] = 16'hFF44;
	assign weights[249] = 16'hFF46;
	assign weights[250] = 16'hFF61;
	assign weights[251] = 16'hFF8C;
	assign weights[252] = 16'hFFBE;
	assign weights[253] = 16'hFFE4;
	assign weights[254] = 16'hFFF5;
	assign weights[255] = 16'hFFED;
endmodule
